module medianSort_N8_k8 ( clk, rst,
dataIn0, dataIn1, dataIn2, dataIn3, dataIn4, dataIn5, dataIn6, dataIn7, dataOut); 

input clk, rst;
input [7:0] dataIn0;
input [7:0] dataIn1;
input [7:0] dataIn2;
input [7:0] dataIn3;
input [7:0] dataIn4;
input [7:0] dataIn5;
input [7:0] dataIn6;
input [7:0] dataIn7;

module medianSort_N16_k8 ( clk, rst,
dataIn0, dataIn1, dataIn2, dataIn3, dataIn4, dataIn5, dataIn6, dataIn7, dataIn8, dataIn9, dataIn10, dataIn11, dataIn12, dataIn13, dataIn14, dataIn15, dataOut); 

input clk, rst;
input [7:0] dataIn0, dataIn1, dataIn2, dataIn3, dataIn4, dataIn5, dataIn6, dataIn7, dataIn8, dataIn9, dataIn10, dataIn11, dataIn12, dataIn13, dataIn14, dataIn15, dataIn16;
